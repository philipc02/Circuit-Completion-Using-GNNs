*SPICE Netlist for circuit 236
I1 1 0 DC 1mA
M4 12 8 1 1 NMOS W=1u L=1u
M3 13 9 1 1 NMOS W=1u L=1u
R2 2 VDD 1k
M1 2 6 12 14 14 NMOS W=1u L=1u
R1 3 VDD 1k
M2 3 6 13 13 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

