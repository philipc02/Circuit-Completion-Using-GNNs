*SPICE Netlist for circuit 755
M6 4 3 0 0 NMOS W=1u L=1u
M3 10 6 0 0 NMOS W=1u L=1u
M7 11 6 0 0 NMOS W=1u L=1u
M8 19 1 VDD 20 20 PMOS W=1u L=1u
M1 9 2 21 22 22 NMOS W=1u L=1u
M5 21 18 4 4 NMOS W=1u L=1u
M2 23 16 4 4 NMOS W=1u L=1u
M10 9 5 19 19 PMOS W=1u L=1u
M13 12 5 24 24 PMOS W=1u L=1u
R2 10 6 1k
R1 6 11 1k
M9 10 9 VDD VDD PMOS W=1u L=1u
M12 11 12 VDD VDD PMOS W=1u L=1u
M4 12 2 23 23 NMOS W=1u L=1u
M11 24 1 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

