*SPICE Netlist for circuit 598
C1 0 2 1nF
M1 1 2 0 0 NMOS W=1u L=1u
R3 0 5 1k
R4 5 1 1k
R2 1 VDD 1k
M2 2 7 5 5 NMOS W=1u L=1u
R1 2 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

