*SPICE Netlist for circuit 631
I1 VDD 1 DC 1mA
I2 2 0 DC 1mA
M1 4 1 8 8 NMOS W=1u L=1u
M3 5 1 9 9 NMOS W=1u L=1u
M5 8 6 2 2 NMOS W=1u L=1u
M2 9 7 2 2 NMOS W=1u L=1u
M4 1 1 2 2 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

