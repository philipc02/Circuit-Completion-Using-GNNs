*SPICE Netlist for circuit 727
C1 1 VDD 1nF
C2 0 3 1nF
C3 10 3 1nF
R2 1 10 1k
M1 6 5 0 12 12 NMOS W=1u L=1u
M2 5 5 0 0 NMOS W=1u L=1u
M3 3 5 0 0 NMOS W=1u L=1u
M5 3 1 VDD VDD PMOS W=1u L=1u
M4 5 6 VDD VDD PMOS W=1u L=1u
M6 6 6 13 13 PMOS W=1u L=1u
R1 13 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

