*SPICE Netlist for circuit 0
M1 1 2 0 0 NMOS W=1u L=1u
V1 2 0 5V
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

