*SPICE Netlist for circuit 219
C1 0 13 1nF
I1 12 0 DC 1mA
I2 3 0 DC 1mA
R1 1 VDD 1k
M4 1 15 3 3 NMOS W=1u L=1u
R2 2 VDD 1k
M3 2 4 14 14 NMOS W=1u L=1u
M2 4 16 3 3 NMOS W=1u L=1u
R3 4 VDD 1k
R4 5 VDD 1k
M1 5 12 8 8 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

