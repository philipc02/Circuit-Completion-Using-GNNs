*SPICE Netlist for circuit 256
R1 0 2 1k
M1 1 4 0 0 NMOS W=1u L=1u
M2 1 1 VDD VDD PMOS W=1u L=1u
M3 2 5 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

