*SPICE Netlist for circuit 276
M3 3 1 0 0 NMOS W=1u L=1u
M4 2 2 VDD VDD NMOS W=1u L=1u
M5 4 2 VDD VDD PMOS W=1u L=1u
M2 2 8 3 3 NMOS W=1u L=1u
M1 4 7 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

