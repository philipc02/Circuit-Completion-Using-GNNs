*SPICE Netlist for circuit 192
M3 1 2 0 0 NMOS W=1u L=1u
M2 6 3 1 1 NMOS W=1u L=1u
M1 7 4 1 1 NMOS W=1u L=1u
R2 7 VDD 1k
R1 6 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

