*SPICE Netlist for circuit 526
I1 2 0 DC 1mA
M3 1 1 VDD VDD NMOS W=1u L=1u
M4 4 1 VDD VDD PMOS W=1u L=1u
M2 1 6 2 2 NMOS W=1u L=1u
M1 4 7 2 2 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

