*SPICE Netlist for circuit 581
I1 0 3 DC 1mA
M1 1 3 0 0 NMOS W=1u L=1u
R2 0 3 1k
R3 3 1 1k
R1 1 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

