*SPICE Netlist for circuit 696
I1 1 0 DC 1mA
M2 2 4 VDD VDD PMOS W=1u L=1u
M1 2 3 1 1 NMOS W=1u L=1u
M3 5 6 2 2 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

