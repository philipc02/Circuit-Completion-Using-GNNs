*SPICE Netlist for circuit 25
M1 4 1 5 5 NMOS W=1u L=1u
V1 4 0 5V
V2 5 0 5V
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

