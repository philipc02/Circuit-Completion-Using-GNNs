*SPICE Netlist for circuit 364
C1 0 3 1nF
C2 0 2 1nF
C3 2 3 1nF
I1 VDD 3 DC 1mA
M1 3 2 0 0 NMOS W=1u L=1u
V1 5 0 5V
R1 5 2 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

