*SPICE Netlist for circuit 265
I1 VDD 2 DC 1mA
M3 6 3 0 0 NMOS W=1u L=1u
M4 1 1 0 0 NMOS W=1u L=1u
M2 4 2 1 1 NMOS W=1u L=1u
R1 4 2 1k
M1 3 4 6 6 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

