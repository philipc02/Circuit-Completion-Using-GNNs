*SPICE Netlist for circuit 735
C1 0 3 1nF
C2 5 3 1nF
I1 4 0 DC 1mA
I2 5 0 DC 1mA
M3 3 4 VDD VDD PMOS W=1u L=1u
M1 3 5 0 0 NMOS W=1u L=1u
M2 4 4 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

