*SPICE Netlist for circuit 140
R1 1 VDD 1k
M1 1 2 5 5 NMOS W=1u L=1u
M2 5 4 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

