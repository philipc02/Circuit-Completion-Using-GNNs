*SPICE Netlist for circuit 416
I1 VDD 3 DC 1mA
I2 1 0 DC 1mA
R1 5 1 1k
M2 3 2 1 1 NMOS W=1u L=1u
M1 VDD 3 1 1 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

