*SPICE Netlist for circuit 813
I1 1 0 DC 1mA
M2 4 7 1 1 NMOS W=1u L=1u
M1 3 8 1 1 NMOS W=1u L=1u
M3 4 2 VDD 10 10 PMOS W=1u L=1u
M4 3 2 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

