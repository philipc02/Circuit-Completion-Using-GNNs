*SPICE Netlist for circuit 56
C1 3 1 1nF
C2 3 2 1nF
V1 2 0 5V
M1 1 3 2 2 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

