*SPICE Netlist for circuit 673
I1 VDD 14 DC 1mA
M6 14 14 0 0 NMOS W=1u L=1u
M7 26 23 0 0 NMOS W=1u L=1u
M3 27 23 0 28 28 NMOS W=1u L=1u
M13 29 1 0 0 NMOS W=1u L=1u
M14 8 12 0 0 NMOS W=1u L=1u
M8 8 11 0 0 NMOS W=1u L=1u
M10 9 5 2 2 NMOS W=1u L=1u
M5 10 6 2 2 NMOS W=1u L=1u
M17 3 3 VDD VDD PMOS W=1u L=1u
M15 9 3 VDD 30 30 PMOS W=1u L=1u
M9 3 6 31 31 NMOS W=1u L=1u
M4 3 18 19 19 NMOS W=1u L=1u
M2 31 32 29 14 14 NMOS W=1u L=1u
M12 2 32 8 8 NMOS W=1u L=1u
M19 12 24 10 10 PMOS W=1u L=1u
M18 10 3 VDD VDD PMOS W=1u L=1u
M16 11 24 9 33 33 PMOS W=1u L=1u
M11 12 25 27 27 NMOS W=1u L=1u
M1 11 25 26 34 34 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

