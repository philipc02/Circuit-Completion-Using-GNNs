*SPICE Netlist for circuit 426
C1 5 VDD 1nF
C2 4 VDD 1nF
I1 1 0 DC 1mA
M2 2 8 1 1 NMOS W=1u L=1u
M1 3 9 1 1 NMOS W=1u L=1u
R2 5 2 1k
M4 2 5 VDD VDD PMOS W=1u L=1u
R1 3 4 1k
M3 3 4 VDD VDD NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

