*SPICE Netlist for circuit 272
I1 2 0 DC 1mA
M1 1 0 2 2 NMOS W=1u L=1u
R1 1 VDD 1k
M2 VDD 4 2 2 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

