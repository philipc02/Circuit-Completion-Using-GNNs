*SPICE Netlist for circuit 730
C1 5 4 1nF
I1 5 0 DC 1mA
I2 3 0 DC 1mA
M5 5 4 VDD VDD PMOS W=1u L=1u
M3 4 2 VDD VDD PMOS W=1u L=1u
M4 2 2 VDD VDD PMOS W=1u L=1u
M2 4 9 3 3 NMOS W=1u L=1u
M1 2 5 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

