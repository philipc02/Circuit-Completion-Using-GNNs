*SPICE Netlist for circuit 618
M1 1 3 0 0 NMOS W=1u L=1u
R3 0 5 1k
R4 3 1 1k
R2 1 VDD 1k
R5 5 1 1k
R1 3 VDD 1k
M2 3 7 5 5 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

