*SPICE Netlist for circuit 307
C1 10 VDD 1nF
C2 8 1 1nF
I1 VDD 2 DC 1mA
I2 3 0 DC 1mA
M2 4 1 0 0 NMOS W=1u L=1u
M1 2 2 0 0 NMOS W=1u L=1u
R1 2 1 1k
R2 3 4 1k
M3 4 10 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

