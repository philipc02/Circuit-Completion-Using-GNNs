*SPICE Netlist for circuit 44
C1 0 1 1nF
I1 4 0 DC 1mA
M1 1 2 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

