*SPICE Netlist for circuit 154
M2 3 1 VDD VDD PMOS W=1u L=1u
M1 3 2 6 6 NMOS W=1u L=1u
R1 5 6 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

