*SPICE Netlist for circuit 718
C1 0 3 1nF
C2 0 5 1nF
I1 4 0 DC 1mA
I2 3 0 DC 1mA
M1 5 3 4 4 NMOS W=1u L=1u
M2 VDD 5 3 3 NMOS W=1u L=1u
M4 2 2 VDD VDD PMOS W=1u L=1u
M5 5 2 VDD VDD PMOS W=1u L=1u
M3 2 8 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

