*SPICE Netlist for circuit 21
C1 7 3 1nF
C2 9 3 1nF
C3 9 7 1nF
C4 9 6 1nF
C5 3 6 1nF
I1 15 7 DC 1mA
I2 6 7 DC 1mA
R1 7 6 1k

.OP
.END

