*SPICE Netlist for circuit 234
I1 2 0 DC 1mA
M1 6 10 1 19 19 NMOS W=1u L=1u
M6 1 12 2 2 NMOS W=1u L=1u
M4 5 13 2 2 NMOS W=1u L=1u
R2 3 VDD 1k
M2 3 11 1 20 20 NMOS W=1u L=1u
M5 3 10 5 5 NMOS W=1u L=1u
M3 6 11 5 5 NMOS W=1u L=1u
R1 6 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

