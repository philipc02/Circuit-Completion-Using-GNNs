*SPICE Netlist for circuit 671
I1 VDD 9 DC 1mA
M5 19 15 0 0 NMOS W=1u L=1u
M2 20 15 0 21 21 NMOS W=1u L=1u
M10 22 1 0 0 NMOS W=1u L=1u
M11 4 8 0 0 NMOS W=1u L=1u
M6 4 7 0 0 NMOS W=1u L=1u
M7 5 10 2 2 NMOS W=1u L=1u
M3 6 11 2 2 NMOS W=1u L=1u
M4 9 9 22 22 NMOS W=1u L=1u
M9 2 9 4 4 NMOS W=1u L=1u
M12 5 16 VDD 23 23 PMOS W=1u L=1u
M14 6 16 VDD VDD PMOS W=1u L=1u
M15 8 17 6 6 PMOS W=1u L=1u
M13 7 17 5 24 24 PMOS W=1u L=1u
M8 8 18 20 20 NMOS W=1u L=1u
M1 7 18 19 25 25 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

