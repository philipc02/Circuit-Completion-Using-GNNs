*SPICE Netlist for circuit 247
I1 1 0 DC 1mA
R3 8 1 1k
R4 1 9 1k
R2 2 VDD 1k
M1 2 5 9 9 NMOS W=1u L=1u
R1 3 VDD 1k
M2 3 7 8 8 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

