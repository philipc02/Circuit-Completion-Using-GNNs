*SPICE Netlist for circuit 394
C1 1 VDD 1nF
C2 0 3 1nF
C3 3 1 1nF
R2 0 3 1k
M1 1 7 0 0 NMOS W=1u L=1u
R1 1 VDD 1k
M2 3 1 VDD VDD PMOS W=1u L=1u
R3 6 7 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

