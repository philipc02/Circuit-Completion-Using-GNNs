*SPICE Netlist for circuit 211
R3 0 2 1k
R1 1 VDD 1k
M1 1 4 2 5 5 NMOS W=1u L=1u
M2 1 4 2 2 NMOS W=1u L=1u
R2 1 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

