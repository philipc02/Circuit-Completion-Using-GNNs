*SPICE Netlist for circuit 280
I1 3 0 DC 1mA
R2 1 3 1k
M4 1 2 VDD VDD PMOS W=1u L=1u
M1 1 8 3 3 NMOS W=1u L=1u
M3 2 2 VDD VDD NMOS W=1u L=1u
M2 2 9 3 3 NMOS W=1u L=1u
R1 3 2 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

