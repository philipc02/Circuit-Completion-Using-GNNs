*SPICE Netlist for circuit 734
C1 0 1 1nF
C2 4 1 1nF
I2 4 0 DC 1mA
I1 VDD 1 DC 1mA

.OP
.END

