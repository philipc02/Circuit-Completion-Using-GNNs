*SPICE Netlist for circuit 1
V1 0 2 5V
M1 1 2 0 0 PMOS W=1u L=1u
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

