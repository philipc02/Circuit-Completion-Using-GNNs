*SPICE Netlist for circuit 642
C1 8 37 1nF
R1 37 1 1k
C2 9 38 1nF
R2 38 2 1k
I1 3 0 DC 1mA
M2 39 34 0 40 40 NMOS W=1u L=1u
M6 41 34 0 0 NMOS W=1u L=1u
R4 6 1 1k
M4 4 1 3 3 NMOS W=1u L=1u
M3 5 2 3 3 NMOS W=1u L=1u
R3 2 7 1k
M8 4 20 VDD VDD PMOS W=1u L=1u
M9 7 35 5 5 PMOS W=1u L=1u
M7 6 35 4 42 42 PMOS W=1u L=1u
M5 7 36 41 41 NMOS W=1u L=1u
M1 6 36 39 43 43 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

