*SPICE Netlist for circuit 753
M5 3 2 0 0 NMOS W=1u L=1u
M1 7 1 13 14 14 NMOS W=1u L=1u
M4 13 12 3 3 NMOS W=1u L=1u
M2 15 10 3 3 NMOS W=1u L=1u
M6 16 4 VDD 17 17 PMOS W=1u L=1u
M7 7 5 16 16 PMOS W=1u L=1u
M9 8 5 18 18 PMOS W=1u L=1u
M3 8 1 15 15 NMOS W=1u L=1u
M8 18 4 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

