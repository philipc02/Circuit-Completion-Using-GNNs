*SPICE Netlist for circuit 32
I1 3 0 DC 1mA
M1 2 1 3 3 NMOS W=1u L=1u
V1 1 0 5V
R1 3 1 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

