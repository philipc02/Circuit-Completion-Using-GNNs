*SPICE Netlist for circuit 181
C1 3 VDD 1nF
M2 4 2 3 3 NMOS W=1u L=1u
M1 VDD 1 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

