*SPICE Netlist for circuit 4
V1 3 0 5V
M1 1 2 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

