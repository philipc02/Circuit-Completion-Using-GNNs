*SPICE Netlist for circuit 785
C1 0 1 1nF
M1 7 3 1 10 10 NMOS W=1u L=1u
M2 2 4 2 2 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

