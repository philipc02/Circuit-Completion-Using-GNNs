*SPICE Netlist for circuit 481
I1 VDD 7 DC 1mA
I2 VDD 4 DC 1mA
I3 4 2 DC 1mA
I4 7 3 DC 1mA
I5 2 0 DC 1mA
M2 4 9 2 2 NMOS W=1u L=1u
M1 7 9 3 3 NMOS W=1u L=1u
R2 7 VDD 1k
R1 4 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

