*SPICE Netlist for circuit 606
V1 4 0 5V
R1 4 1 1k
R2 1 1 1k

.OP
.END

