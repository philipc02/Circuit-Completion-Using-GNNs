*SPICE Netlist for circuit 77
M2 1 3 0 0 NMOS W=1u L=1u
M1 VDD VDD 1 1 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

