*SPICE Netlist for circuit 134
I1 VDD 2 DC 1mA
M2 5 4 0 0 NMOS W=1u L=1u
M1 2 1 5 5 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

