*SPICE Netlist for circuit 690
C1 5 3 1nF
C2 0 5 1nF
I1 4 0 DC 1mA
M2 1 1 VDD VDD PMOS W=1u L=1u
M3 3 1 VDD VDD PMOS W=1u L=1u
M1 1 8 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

