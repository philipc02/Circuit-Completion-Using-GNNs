*SPICE Netlist for circuit 512
R2 0 4 1k
M2 2 1 VDD VDD PMOS W=1u L=1u
R1 4 2 1k
M1 2 6 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

