*SPICE Netlist for circuit 650
V1 1 0 5V
R2 0 2 1k
R1 2 1 1k

.OP
.END

