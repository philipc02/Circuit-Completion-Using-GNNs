*SPICE Netlist for circuit 94
R3 0 1 1k
R2 0 1 1k
R1 2 1 1k

.OP
.END

