*SPICE Netlist for circuit 39
V1 5 0 5V
V2 4 0 5V
M1 2 1 5 5 NMOS W=1u L=1u
R1 2 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

