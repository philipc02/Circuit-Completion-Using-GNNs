*SPICE Netlist for circuit 657
I1 4 0 DC 1mA
M3 2 1 VDD VDD PMOS W=1u L=1u
M2 2 2 4 4 NMOS W=1u L=1u
M1 3 3 4 4 NMOS W=1u L=1u
M4 3 7 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

