*SPICE Netlist for circuit 8
I1 VDD 1 DC 1mA

.OP
.END

