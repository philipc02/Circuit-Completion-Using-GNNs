*SPICE Netlist for circuit 522
I1 2 0 DC 1mA
M2 1 2 0 0 NMOS W=1u L=1u
M1 VDD 1 2 2 NMOS W=1u L=1u
R1 1 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

