*SPICE Netlist for circuit 180
I1 3 0 DC 1mA
M2 2 5 0 0 NMOS W=1u L=1u
M1 VDD 2 3 3 NMOS W=1u L=1u
M3 2 3 VDD VDD NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

