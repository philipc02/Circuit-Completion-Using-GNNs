*SPICE Netlist for circuit 348
I1 2 0 DC 1mA
M3 1 1 VDD VDD NMOS W=1u L=1u
M4 6 1 VDD VDD PMOS W=1u L=1u
M1 6 8 2 2 NMOS W=1u L=1u
M2 1 9 2 2 NMOS W=1u L=1u
R1 2 1 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

