*SPICE Netlist for circuit 796
C1 0 2 1nF
C2 0 1 1nF
M1 6 3 1 1 NMOS W=1u L=1u
M2 1 4 2 2 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

