*SPICE Netlist for circuit 291
I1 2 0 DC 1mA
I2 3 0 DC 1mA
M1 2 2 VDD VDD NMOS W=1u L=1u
M2 3 2 VDD VDD PMOS W=1u L=1u
R1 2 VDD 1k
R2 3 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

