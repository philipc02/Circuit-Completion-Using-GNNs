*SPICE Netlist for circuit 737
C1 2 1nF
I1 VDD 4 DC 1mA
I2 VDD 2 DC 1mA
I3 3 0 DC 1mA
M1 6 3 0 0 NMOS W=1u L=1u
M3 3 1 4 4 PMOS W=1u L=1u
M2 3 7 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

