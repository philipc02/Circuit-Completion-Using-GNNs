*SPICE Netlist for circuit 193
I1 2 0 DC 1mA
R2 1 VDD 1k
M1 1 5 2 2 NMOS W=1u L=1u
M2 3 7 2 2 NMOS W=1u L=1u
R1 3 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

