*SPICE Netlist for circuit 788
I1 1 0 DC 1mA
V1 4 0 5V
R2 4 1 1k
R1 0 1 1k

.OP
.END

