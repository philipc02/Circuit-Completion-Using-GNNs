*SPICE Netlist for circuit 652
I1 VDD 3 DC 1mA
I2 2 0 DC 1mA
M2 1 5 0 0 NMOS W=1u L=1u
M3 2 1 6 6 PMOS W=1u L=1u
M1 3 2 1 1 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

