*SPICE Netlist for circuit 577
R6 4 0 1k
R2 0 4 1k
R3 0 1 1k
R4 0 2 1k
R5 1 2 1k
M2 2 3 VDD VDD PMOS W=1u L=1u
R1 3 VDD 1k
M1 3 5 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

