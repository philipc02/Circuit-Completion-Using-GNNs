*SPICE Netlist for circuit 245
M3 2 3 0 0 NMOS W=1u L=1u
M4 1 5 VDD VDD PMOS W=1u L=1u
M2 1 12 2 2 NMOS W=1u L=1u
M1 5 10 2 2 NMOS W=1u L=1u
M6 1 1 VDD VDD PMOS W=1u L=1u
M5 5 5 VDD VDD PMOS W=1u L=1u
M7 5 1 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

