*SPICE Netlist for circuit 57
M1 2 1 5 5 NMOS W=1u L=1u
M2 5 1 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

