*SPICE Netlist for circuit 467
I1 VDD 4 DC 1mA
I2 4 3 DC 1mA
M1 4 1 3 3 NMOS W=1u L=1u
R1 4 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

