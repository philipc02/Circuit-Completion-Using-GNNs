*SPICE Netlist for circuit 405
C1 2 5 1nF
C2 0 3 1nF
C3 5 3 1nF
I1 3 2 DC 1mA
R3 0 5 1k
R1 0 3 1k
V1 7 0 5V
R2 7 2 1k

.OP
.END

