*SPICE Netlist for circuit 821
C1 0 3 1nF
C2 0 2 1nF
C3 0 4 1nF
M1 2 4 0 0 NMOS W=1u L=1u
M2 3 2 0 0 NMOS W=1u L=1u
M3 4 3 0 0 NMOS W=1u L=1u
R1 2 VDD 1k
R2 3 VDD 1k
R3 4 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

