*SPICE Netlist for circuit 582
I1 0 2 DC 1mA
R4 0 1 1k
M1 1 2 0 0 NMOS W=1u L=1u
R3 0 2 1k
R2 2 0 1k
R1 1 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

