*SPICE Netlist for circuit 99
I1 1 0 DC 1mA
M1 VDD 3 1 1 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

