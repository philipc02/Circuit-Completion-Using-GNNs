*SPICE Netlist for circuit 164
I1 VDD 3 DC 1mA
V1 6 0 5V
M1 6 1 3 3 NMOS W=1u L=1u
M2 3 2 0 0 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

