*SPICE Netlist for circuit 215
V2 4 0 5V
R3 0 2 1k
R1 1 VDD 1k
M2 1 9 2 2 NMOS W=1u L=1u
M1 3 4 2 2 NMOS W=1u L=1u
R2 3 VDD 1k
V1 9 4 5V
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

