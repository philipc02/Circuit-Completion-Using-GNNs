*SPICE Netlist for circuit 741
C1 0 2 1nF
C2 0 4 1nF
I1 3 0 DC 1mA
I2 4 0 DC 1mA
M4 2 1 VDD VDD PMOS W=1u L=1u
M2 VDD 2 4 4 NMOS W=1u L=1u
M3 VDD 8 3 3 NMOS W=1u L=1u
M1 2 9 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

