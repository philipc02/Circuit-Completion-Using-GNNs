*SPICE Netlist for circuit 358
I1 VDD 2 DC 1mA
R2 3 0 1k
M1 2 1 3 3 NMOS W=1u L=1u
R1 2 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

