*SPICE Netlist for circuit 483
I1 1 2 DC 1mA
R2 1 VDD 1k
R1 0 2 1k
M1 1 3 2 2 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

