*SPICE Netlist for circuit 257
I1 VDD 3 DC 1mA
M3 VDD 3 6 6 NMOS W=1u L=1u
M2 2 2 0 0 NMOS W=1u L=1u
M4 6 2 0 0 NMOS W=1u L=1u
M1 3 3 2 2 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

