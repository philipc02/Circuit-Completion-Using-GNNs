*SPICE Netlist for circuit 769
M1 3 3 0 0 NMOS W=1u L=1u
M2 1 5 0 0 NMOS W=1u L=1u
M3 5 6 0 0 NMOS W=1u L=1u
R1 8 0 1k
M5 3 1 VDD VDD PMOS W=1u L=1u
M6 1 1 VDD VDD PMOS W=1u L=1u
M4 1 3 8 8 NMOS W=1u L=1u
R3 5 6 1k
R2 6 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

