*SPICE Netlist for circuit 450
I1 1 3 DC 1mA
M1 1 5 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

