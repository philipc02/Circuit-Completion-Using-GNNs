*SPICE Netlist for circuit 283
V1 3 0 5V
M1 3 0 5 5 NMOS W=1u L=1u
M2 1 0 5 5 NMOS W=1u L=1u
M3 1 1 VDD VDD NMOS W=1u L=1u
M4 3 1 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

