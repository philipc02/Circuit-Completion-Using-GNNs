*SPICE Netlist for circuit 341
C1 3 1 1nF
M1 1 1 3 3 NMOS W=1u L=1u
M2 4 1 0 0 NMOS W=1u L=1u
R1 1 VDD 1k
R2 4 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

