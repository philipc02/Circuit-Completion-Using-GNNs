*SPICE Netlist for circuit 267
I1 VDD 3 DC 1mA
V1 2 0 5V
M1 3 3 0 0 NMOS W=1u L=1u
M3 2 3 0 0 NMOS W=1u L=1u
M2 3 2 0 0 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

