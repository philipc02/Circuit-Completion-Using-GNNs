*SPICE Netlist for circuit 508
I1 VDD 2 DC 1mA
R2 0 3 1k
R1 3 2 1k
M1 2 5 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

