*SPICE Netlist for circuit 803
C1 0 3 1nF
M2 3 1 5 5 PMOS W=1u L=1u
M1 3 4 5 5 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

