*SPICE Netlist for circuit 35
R1 0 2 1k
V1 4 0 5V
M1 2 1 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

