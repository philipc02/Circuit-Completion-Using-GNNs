*SPICE Netlist for circuit 681
I1 3 0 DC 1mA
M2 8 5 0 0 NMOS W=1u L=1u
M4 9 5 0 0 NMOS W=1u L=1u
M6 8 1 VDD VDD PMOS W=1u L=1u
R4 1 2 1k
M5 1 2 VDD VDD PMOS W=1u L=1u
M3 1 13 3 3 NMOS W=1u L=1u
M7 7 2 VDD VDD PMOS W=1u L=1u
M1 7 14 3 3 NMOS W=1u L=1u
R1 2 7 1k
R2 8 5 1k
R3 5 9 1k
M8 9 7 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

