*SPICE Netlist for circuit 817
I1 1 0 DC 1mA
M4 11 10 1 1 NMOS W=1u L=1u
M2 12 8 1 1 NMOS W=1u L=1u
M1 4 2 11 13 13 NMOS W=1u L=1u
R2 3 VDD 1k
M3 3 2 12 12 NMOS W=1u L=1u
R1 4 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

