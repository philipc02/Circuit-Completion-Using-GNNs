*SPICE Netlist for circuit 60
V1 2 0 5V
M1 2 3 1 5 5 NMOS W=1u L=1u
M2 1 3 2 2 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

