*SPICE Netlist for circuit 384
M3 1 2 0 0 NMOS W=1u L=1u
M2 4 8 1 1 NMOS W=1u L=1u
M1 3 6 1 1 NMOS W=1u L=1u
R2 3 VDD 1k
R1 4 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

