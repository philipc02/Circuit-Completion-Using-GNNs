*SPICE Netlist for circuit 20
M1 3 8 1 1 NMOS W=1u L=1u
M2 3 9 1 1 NMOS W=1u L=1u
R1 5 8 1k
R2 9 5 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

