*SPICE Netlist for circuit 404
C1 2 5 1nF
C2 0 3 1nF
C3 5 3 1nF
I1 3 2 DC 1mA
V1 7 0 5V
R1 0 3 1k
R2 0 2 1k
R3 7 5 1k

.OP
.END

