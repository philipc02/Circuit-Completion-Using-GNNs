*SPICE Netlist for circuit 320
M5 3 1 0 0 NMOS W=1u L=1u
M6 4 2 0 0 NMOS W=1u L=1u
M3 8 11 3 3 NMOS W=1u L=1u
M1 6 12 3 3 NMOS W=1u L=1u
M4 7 6 4 4 NMOS W=1u L=1u
M2 5 8 4 4 NMOS W=1u L=1u
R4 5 VDD 1k
R2 6 VDD 1k
R3 7 VDD 1k
R1 8 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

