*SPICE Netlist for circuit 472
C1 0 6 1nF
C2 0 1 1nF
I1 VDD 1 DC 1mA
I2 6 0 DC 1mA
I3 3 0 DC 1mA
M2 3 1 0 0 NMOS W=1u L=1u
M3 1 1 0 0 NMOS W=1u L=1u
M1 4 5 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

