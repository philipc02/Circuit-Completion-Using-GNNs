*SPICE Netlist for circuit 299
C1 5 2 1nF
M1 3 2 0 0 NMOS W=1u L=1u
R2 1 2 1k
R1 3 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

