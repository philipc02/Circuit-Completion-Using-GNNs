*SPICE Netlist for circuit 255
I1 VDD 7 DC 1mA
M3 7 7 0 0 NMOS W=1u L=1u
M1 1 7 0 8 8 NMOS W=1u L=1u
M5 1 1 VDD VDD NMOS W=1u L=1u
M8 3 1 VDD VDD PMOS W=1u L=1u
M9 2 2 VDD VDD PMOS W=1u L=1u
M7 2 VDD VDD VDD NMOS W=1u L=1u
M2 2 9 4 4 NMOS W=1u L=1u
M6 3 3 VDD VDD NMOS W=1u L=1u
M4 3 10 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

