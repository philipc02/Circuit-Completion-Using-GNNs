*SPICE Netlist for circuit 121
I1 VDD 3 DC 1mA
V1 6 0 5V
M1 3 1 4 4 NMOS W=1u L=1u
R2 4 3 1k
R1 6 4 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

