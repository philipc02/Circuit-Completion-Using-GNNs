*SPICE Netlist for circuit 596
M1 2 1 0 0 NMOS W=1u L=1u
M2 1 0 4 4 NMOS W=1u L=1u
R1 0 4 1k
V1 7 0 5V
R3 1 VDD 1k
R2 2 VDD 1k
R4 4 7 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

