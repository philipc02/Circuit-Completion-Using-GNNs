*SPICE Netlist for circuit 295
I1 3 0 DC 1mA
V1 2 0 5V
M3 1 1 VDD VDD NMOS W=1u L=1u
M4 5 1 VDD VDD PMOS W=1u L=1u
M2 1 2 3 3 NMOS W=1u L=1u
M1 5 2 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

