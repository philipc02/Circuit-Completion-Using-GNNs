*SPICE Netlist for circuit 521
M1 2 3 0 0 NMOS W=1u L=1u
R1 0 3 1k
M2 3 1 2 2 PMOS W=1u L=1u
R2 2 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

