*SPICE Netlist for circuit 58


.OP
.END

