*SPICE Netlist for circuit 395
C1 3 VDD 1nF
C2 0 1 1nF
R2 0 1 1k
M1 3 6 0 0 NMOS W=1u L=1u
M2 1 3 VDD VDD PMOS W=1u L=1u
R1 3 VDD 1k
R3 5 6 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

