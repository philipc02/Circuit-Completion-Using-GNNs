*SPICE Netlist for circuit 432
I1 1 4 DC 1mA
I2 3 6 DC 1mA
R1 1 4 1k
R2 4 1 1k

.OP
.END

