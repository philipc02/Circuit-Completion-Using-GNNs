*SPICE Netlist for circuit 651
I1 VDD 3 DC 1mA
I2 VDD 2 DC 1mA
M1 3 1 0 0 NMOS W=1u L=1u
M3 1 5 0 0 NMOS W=1u L=1u
M2 2 3 1 1 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

