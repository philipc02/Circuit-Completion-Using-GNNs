*SPICE Netlist for circuit 716
I1 VDD 5 DC 1mA
M2 4 22 0 0 NMOS W=1u L=1u
M4 2 20 0 0 NMOS W=1u L=1u
M3 7 3 0 0 NMOS W=1u L=1u
M5 11 8 0 0 NMOS W=1u L=1u
M1 3 1 0 23 23 NMOS W=1u L=1u
M6 8 1 0 0 NMOS W=1u L=1u
M8 2 2 VDD VDD PMOS W=1u L=1u
M11 11 2 VDD VDD PMOS W=1u L=1u
M7 7 4 VDD VDD PMOS W=1u L=1u
M10 4 4 VDD VDD PMOS W=1u L=1u
M12 3 15 5 5 PMOS W=1u L=1u
M9 8 16 5 5 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

