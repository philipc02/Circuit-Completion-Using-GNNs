*SPICE Netlist for circuit 608
I1 VDD 2 DC 1mA
I2 1 0 DC 1mA
M2 2 1 0 0 NMOS W=1u L=1u
R1 4 1 1k
M1 VDD 2 1 1 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

