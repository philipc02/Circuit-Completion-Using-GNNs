*SPICE Netlist for circuit 764
V1 VDD 0 5V
R4 0 3 1k
R5 0 6 1k
M2 3 1 2 2 NMOS W=1u L=1u
R1 1 VDD 1k
R2 2 3 1k
R3 6 1 1k
M1 1 3 6 6 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

