*SPICE Netlist for circuit 117
V1 2 0 5V
R1 2 1 1k

.OP
.END

