*SPICE Netlist for circuit 198
R1 0 4 1k
R2 1 VDD 1k
M1 1 3 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

