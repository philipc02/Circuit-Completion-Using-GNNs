*SPICE Netlist for circuit 635
I1 VDD 2 DC 1mA
I2 3 0 DC 1mA
M1 2 5 0 0 NMOS W=1u L=1u
M2 3 1 2 2 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

