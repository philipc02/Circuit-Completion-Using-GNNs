*SPICE Netlist for circuit 138
M2 5 1 2 2 NMOS W=1u L=1u
M1 4 1 5 5 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

