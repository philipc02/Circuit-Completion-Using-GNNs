*SPICE Netlist for circuit 469
I1 VDD 3 DC 1mA
I2 7 1 DC 1mA
M1 14 2 1 1 NMOS W=1u L=1u
R1 4 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

