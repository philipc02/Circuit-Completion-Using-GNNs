*SPICE Netlist for circuit 434
I1 VDD 2 DC 1mA
I2 2 3 DC 1mA
M1 2 0 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

