*SPICE Netlist for circuit 459
I1 VDD 2 DC 1mA
I2 2 0 DC 1mA
M1 2 6 0 0 NMOS W=1u L=1u
R1 0 2 1k
M2 2 1 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

