*SPICE Netlist for circuit 298
M1 3 1 0 0 NMOS W=1u L=1u
R1 3 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

