*SPICE Netlist for circuit 23
C1 0 1 1nF
M1 1 2 VDD VDD PMOS W=1u L=1u
V1 VDD 2 5V
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

