*SPICE Netlist for circuit 421
C1 5 1 1nF
I1 3 0 DC 1mA
M4 1 2 VDD VDD PMOS W=1u L=1u
M1 1 8 3 3 NMOS W=1u L=1u
M3 5 2 VDD VDD NMOS W=1u L=1u
M2 5 7 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

