*SPICE Netlist for circuit 195
I1 2 0 DC 1mA
V2 6 0 5V
V1 7 0 5V
R2 1 VDD 1k
M1 1 7 2 2 NMOS W=1u L=1u
M2 3 6 2 2 NMOS W=1u L=1u
R1 3 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

