*SPICE Netlist for circuit 410
I1 VDD 3 DC 1mA
I2 VDD 1 DC 1mA
M2 1 3 0 0 NMOS W=1u L=1u
M1 3 2 6 6 NMOS W=1u L=1u
R1 5 6 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

