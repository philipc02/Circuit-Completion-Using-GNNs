*SPICE Netlist for circuit 253
M1 1 5 0 0 NMOS W=1u L=1u
M3 1 1 VDD VDD PMOS W=1u L=1u
M2 1 3 VDD VDD NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

