*SPICE Netlist for circuit 683
I1 1 0 DC 1mA
M2 13 5 0 14 14 NMOS W=1u L=1u
M6 15 5 0 0 NMOS W=1u L=1u
M4 2 7 1 1 NMOS W=1u L=1u
M3 3 4 1 1 NMOS W=1u L=1u
M8 2 16 VDD VDD PMOS W=1u L=1u
M9 3 10 16 16 PMOS W=1u L=1u
M10 4 12 3 3 PMOS W=1u L=1u
M5 4 11 15 15 NMOS W=1u L=1u
M1 5 11 13 17 17 NMOS W=1u L=1u
M7 5 12 2 18 18 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

