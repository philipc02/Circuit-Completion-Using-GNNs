*SPICE Netlist for circuit 669
M6 17 13 0 0 NMOS W=1u L=1u
M3 18 13 0 19 19 NMOS W=1u L=1u
M10 3 7 0 0 NMOS W=1u L=1u
M7 3 6 0 0 NMOS W=1u L=1u
M8 4 8 1 1 NMOS W=1u L=1u
M4 5 9 1 1 NMOS W=1u L=1u
M5 1 2 3 3 NMOS W=1u L=1u
M12 4 14 VDD VDD PMOS W=1u L=1u
M2 5 14 VDD 20 20 NMOS W=1u L=1u
M13 7 15 5 5 PMOS W=1u L=1u
M11 6 15 4 21 21 PMOS W=1u L=1u
M9 7 16 18 18 NMOS W=1u L=1u
M1 6 16 17 22 22 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

