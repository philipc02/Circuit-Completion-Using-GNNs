*SPICE Netlist for circuit 337
C1 0 3 1nF
M1 2 2 3 3 NMOS W=1u L=1u
I1 VDD 2 DC 1mA
M2 4 2 0 0 NMOS W=1u L=1u
R1 4 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

