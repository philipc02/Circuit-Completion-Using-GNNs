*SPICE Netlist for circuit 225
I1 1 0 DC 1mA
M4 4 2 VDD VDD PMOS W=1u L=1u
M3 6 3 VDD VDD PMOS W=1u L=1u
M2 4 10 1 1 NMOS W=1u L=1u
M1 6 11 1 1 NMOS W=1u L=1u
R1 4 VDD 1k
R2 6 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

