*SPICE Netlist for circuit 104
M2 1 2 0 0 NMOS W=1u L=1u
R1 0 1 1k
M1 VDD 5 1 1 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

