*SPICE Netlist for circuit 353
C1 2 5 1nF
I1 2 0 DC 1mA
M2 3 1 2 2 NMOS W=1u L=1u
M1 5 1 2 2 NMOS W=1u L=1u
M3 3 3 VDD VDD NMOS W=1u L=1u
M4 5 3 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

