*SPICE Netlist for circuit 659
I1 VDD 2 DC 1mA
I2 2 0 DC 1mA
R2 0 2 1k
R1 2 VDD 1k

.OP
.END

