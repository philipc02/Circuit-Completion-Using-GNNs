*SPICE Netlist for circuit 114
V1 6 0 5V
M1 2 1 4 4 NMOS W=1u L=1u
R1 2 VDD 1k
R2 4 2 1k
R3 6 4 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

