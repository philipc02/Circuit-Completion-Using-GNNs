*SPICE Netlist for circuit 324
M2 3 1 0 0 NMOS W=1u L=1u
R1 0 4 1k
M1 1 1 4 4 NMOS W=1u L=1u
R2 1 VDD 1k
R3 3 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

