*SPICE Netlist for circuit 768
M2 2 4 0 0 NMOS W=1u L=1u
M1 4 3 0 0 NMOS W=1u L=1u
M3 3 2 VDD VDD PMOS W=1u L=1u
M4 2 2 VDD VDD PMOS W=1u L=1u
R1 4 3 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

