*SPICE Netlist for circuit 28
M1 2 1 5 5 NMOS W=1u L=1u
V2 5 0 5V
V1 3 0 5V
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

