*SPICE Netlist for circuit 723
C1 1 VDD 1nF
C2 0 3 1nF
R2 0 1 1k
R1 0 1 1k
M1 1 1 VDD VDD PMOS W=1u L=1u
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

