*SPICE Netlist for circuit 48
C1 0 3 1nF
C2 3 2 1nF
M1 2 1 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

