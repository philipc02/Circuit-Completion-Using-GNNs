*SPICE Netlist for circuit 206
I1 2 0 DC 1mA
V1 8 0 5V
V2 9 0 5V
R4 1 2 1k
R2 1 VDD 1k
M1 1 9 2 2 NMOS W=1u L=1u
R3 2 3 1k
R1 3 VDD 1k
M2 3 8 2 2 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

