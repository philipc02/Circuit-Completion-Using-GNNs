*SPICE Netlist for circuit 122
I1 VDD 1 DC 1mA
V1 4 0 5V
M1 1 2 4 4 NMOS W=1u L=1u
R1 4 1 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

