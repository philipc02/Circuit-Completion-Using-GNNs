*SPICE Netlist for circuit 373
C1 1 3 1nF
C2 3 4 1nF
R1 2 4 1k

.OP
.END

