*SPICE Netlist for circuit 686
C1 0 5 1nF
I1 4 0 DC 1mA
M4 2 7 VDD VDD PMOS W=1u L=1u
M2 7 9 4 4 NMOS W=1u L=1u
M1 2 6 4 4 NMOS W=1u L=1u
R1 0 6 1k
M3 7 7 VDD VDD PMOS W=1u L=1u
R2 6 5 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

