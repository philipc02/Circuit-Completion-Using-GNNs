*SPICE Netlist for circuit 106
M2 0 4 2 2 PMOS W=1u L=1u
M1 2 1 VDD VDD PMOS W=1u L=1u
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

