*SPICE Netlist for circuit 150
R1 0 1 1k
R2 2 1 1k
M1 VDD 2 1 1 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

