*SPICE Netlist for circuit 65
R2 0 1 1k
R1 1 VDD 1k

.OP
.END

