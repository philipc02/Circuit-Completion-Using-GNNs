*SPICE Netlist for circuit 519
R3 0 2 1k
R2 2 1 1k
M1 1 2 5 5 NMOS W=1u L=1u
R1 1 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

