*SPICE Netlist for circuit 762
M3 4 3 VDD VDD NMOS W=1u L=1u
M2 3 4 7 7 NMOS W=1u L=1u
M1 4 4 0 0 NMOS W=1u L=1u
R1 0 7 1k
M4 3 3 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

