*SPICE Netlist for circuit 516
R2 5 1 1k
R1 2 VDD 1k
M1 2 5 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

