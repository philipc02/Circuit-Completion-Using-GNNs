*SPICE Netlist for circuit 365
C1 0 2 1nF
C2 2 1 1nF
V1 4 0 5V
M1 1 2 0 0 NMOS W=1u L=1u
R1 1 VDD 1k
R2 4 2 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

