*SPICE Netlist for circuit 676
I1 6 0 DC 1mA
M4 3 5 0 0 NMOS W=1u L=1u
M2 3 2 0 0 NMOS W=1u L=1u
M6 6 6 VDD VDD PMOS W=1u L=1u
M5 5 6 VDD 9 9 PMOS W=1u L=1u
M7 2 6 VDD VDD PMOS W=1u L=1u
M1 2 7 3 3 NMOS W=1u L=1u
M3 5 8 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

