*SPICE Netlist for circuit 643
I1 5 0 DC 1mA
M1 4 1 12 13 13 NMOS W=1u L=1u
M5 2 2 VDD VDD PMOS W=1u L=1u
M6 4 4 2 2 PMOS W=1u L=1u
M7 14 2 VDD VDD PMOS W=1u L=1u
M8 6 4 14 14 PMOS W=1u L=1u
M4 12 9 5 5 NMOS W=1u L=1u
M2 15 10 5 5 NMOS W=1u L=1u
M3 6 1 15 15 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

