*SPICE Netlist for circuit 712
I1 4 0 DC 1mA
M1 5 1 0 12 12 NMOS W=1u L=1u
M4 6 1 0 0 NMOS W=1u L=1u
M6 5 2 VDD VDD PMOS W=1u L=1u
M5 2 2 VDD VDD PMOS W=1u L=1u
M3 2 8 4 4 NMOS W=1u L=1u
M7 3 3 VDD VDD PMOS W=1u L=1u
M8 6 3 VDD VDD PMOS W=1u L=1u
M2 3 9 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

