*SPICE Netlist for circuit 682
I1 9 0 DC 1mA
M7 7 4 0 0 NMOS W=1u L=1u
M3 7 5 0 0 NMOS W=1u L=1u
M4 13 9 0 0 NMOS W=1u L=1u
M8 14 9 0 0 NMOS W=1u L=1u
M9 4 2 VDD 23 23 PMOS W=1u L=1u
M1 4 3 24 25 25 NMOS W=1u L=1u
M10 13 4 VDD VDD PMOS W=1u L=1u
M11 5 2 VDD VDD PMOS W=1u L=1u
M5 5 3 26 26 NMOS W=1u L=1u
M12 14 5 VDD VDD PMOS W=1u L=1u
M6 24 21 7 7 NMOS W=1u L=1u
M2 26 22 7 7 NMOS W=1u L=1u
R1 13 9 1k
R2 9 14 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

