*SPICE Netlist for circuit 300
C1 6 1 1nF
I1 VDD 2 DC 1mA
M2 4 1 0 0 NMOS W=1u L=1u
M1 2 2 0 0 NMOS W=1u L=1u
R2 2 1 1k
R1 4 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

