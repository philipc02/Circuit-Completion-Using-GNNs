*SPICE Netlist for circuit 609
I1 VDD 1 DC 1mA
I2 3 0 DC 1mA
M1 1 3 0 0 NMOS W=1u L=1u
M2 3 2 1 1 PMOS W=1u L=1u
R1 5 3 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

