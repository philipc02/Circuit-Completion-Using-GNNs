*SPICE Netlist for circuit 418
C1 5 4 1nF
M2 5 7 0 0 NMOS W=1u L=1u
M3 4 1 VDD VDD PMOS W=1u L=1u
M1 4 2 5 5 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

