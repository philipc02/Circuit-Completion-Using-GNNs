*SPICE Netlist for circuit 414
I1 VDD 1 DC 1mA
I2 2 0 DC 1mA
M2 2 1 VDD VDD PMOS W=1u L=1u
M1 1 3 2 2 NMOS W=1u L=1u
R1 5 2 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

