*SPICE Netlist for circuit 645
I1 4 0 DC 1mA
M1 6 1 0 14 14 NMOS W=1u L=1u
M4 8 1 0 0 NMOS W=1u L=1u
M5 5 2 VDD VDD NMOS W=1u L=1u
M7 7 2 VDD VDD PMOS W=1u L=1u
M3 5 10 4 4 NMOS W=1u L=1u
M2 7 11 4 4 NMOS W=1u L=1u
M6 6 5 VDD VDD NMOS W=1u L=1u
M8 8 7 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

