*SPICE Netlist for circuit 784
C1 0 1 1nF
R1 3 1 1k

.OP
.END

