*SPICE Netlist for circuit 592
R2 0 1 1k
M1 VDD 2 1 1 NMOS W=1u L=1u
R1 2 VDD 1k
M2 2 5 1 1 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

