*SPICE Netlist for circuit 602
R2 0 1 1k
M1 2 1 0 0 NMOS W=1u L=1u
R3 1 4 1k
V1 3 2 5V
R1 2 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

