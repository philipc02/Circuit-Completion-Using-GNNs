*SPICE Netlist for circuit 216
C1 0 10 1nF
I1 9 0 DC 1mA
M2 2 1 11 11 NMOS W=1u L=1u
R1 2 VDD 1k
R2 3 VDD 1k
M1 3 9 7 7 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

