*SPICE Netlist for circuit 591
M1 2 1 3 3 NMOS W=1u L=1u
R2 3 2 1k
R1 2 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

