*SPICE Netlist for circuit 617
M1 2 5 0 0 NMOS W=1u L=1u
R2 0 3 1k
M3 5 1 VDD 8 8 PMOS W=1u L=1u
R1 3 2 1k
M2 5 7 3 3 NMOS W=1u L=1u
M4 2 1 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

