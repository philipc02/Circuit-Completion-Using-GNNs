*SPICE Netlist for circuit 684
I1 1 0 DC 1mA
M2 8 6 0 21 21 NMOS W=1u L=1u
M7 7 6 0 0 NMOS W=1u L=1u
M5 3 5 1 1 NMOS W=1u L=1u
M4 4 9 1 1 NMOS W=1u L=1u
M12 8 5 2 2 PMOS W=1u L=1u
M10 16 9 2 2 PMOS W=1u L=1u
M9 3 18 VDD VDD PMOS W=1u L=1u
M3 4 18 VDD 22 22 NMOS W=1u L=1u
M11 10 19 4 4 PMOS W=1u L=1u
M8 6 19 3 23 23 PMOS W=1u L=1u
M1 6 20 7 24 24 NMOS W=1u L=1u
M6 10 20 7 7 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

