*SPICE Netlist for circuit 243
M1 8 2 0 14 14 NMOS W=1u L=1u
M4 7 2 0 0 NMOS W=1u L=1u
M6 4 1 VDD VDD PMOS W=1u L=1u
M2 5 3 8 15 15 NMOS W=1u L=1u
M7 8 12 4 4 PMOS W=1u L=1u
M5 7 10 4 4 PMOS W=1u L=1u
R2 5 VDD 1k
R1 6 VDD 1k
M3 6 3 7 7 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

