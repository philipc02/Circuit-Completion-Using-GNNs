*SPICE Netlist for circuit 387
C1 0 1 1nF
C2 2 0 1nF
I1 5 0 DC 1mA
I2 4 0 DC 1mA
M3 1 5 VDD 11 11 PMOS W=1u L=1u
M2 1 8 4 4 NMOS W=1u L=1u
M5 2 5 VDD VDD PMOS W=1u L=1u
M1 2 9 4 4 NMOS W=1u L=1u
M4 5 5 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

