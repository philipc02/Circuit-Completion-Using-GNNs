*SPICE Netlist for circuit 179
M2 2 5 0 0 NMOS W=1u L=1u
M1 6 1 2 2 NMOS W=1u L=1u
M3 6 2 VDD VDD NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

