*SPICE Netlist for circuit 524
I1 1 0 DC 1mA
M1 2 1 0 0 NMOS W=1u L=1u
M2 VDD 2 1 1 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

