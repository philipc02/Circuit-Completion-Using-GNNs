*SPICE Netlist for circuit 230
M2 3 6 1 1 NMOS W=1u L=1u
M1 2 7 1 1 NMOS W=1u L=1u
R2 2 VDD 1k
R1 3 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

