*SPICE Netlist for circuit 232
I1 3 0 DC 1mA
M4 4 11 1 1 NMOS W=1u L=1u
M1 5 13 1 1 NMOS W=1u L=1u
M5 5 12 2 2 NMOS W=1u L=1u
M2 7 14 2 2 NMOS W=1u L=1u
M6 1 15 3 3 NMOS W=1u L=1u
M3 2 10 3 3 NMOS W=1u L=1u
R1 4 VDD 1k
R2 7 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

