*SPICE Netlist for circuit 710
M7 4 3 0 0 NMOS W=1u L=1u
M4 18 6 0 0 NMOS W=1u L=1u
M2 19 6 0 20 20 NMOS W=1u L=1u
V1 17 0 5V
M8 10 1 7 21 21 PMOS W=1u L=1u
M1 10 2 18 22 22 NMOS W=1u L=1u
M5 7 13 4 4 NMOS W=1u L=1u
M3 8 14 4 4 NMOS W=1u L=1u
M10 8 5 VDD VDD PMOS W=1u L=1u
M9 7 23 VDD VDD PMOS W=1u L=1u
M11 9 1 8 8 PMOS W=1u L=1u
M6 9 2 19 19 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

