*SPICE Netlist for circuit 739
C1 0 1 1nF
C2 4 1 1nF
I1 0 4 DC 1mA
R2 0 1 1k
R1 3 0 1k
M2 1 3 0 0 PMOS W=1u L=1u
M1 3 0 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

