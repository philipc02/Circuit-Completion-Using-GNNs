*SPICE Netlist for circuit 235
I1 1 0 DC 1mA
M4 11 8 1 1 NMOS W=1u L=1u
M2 12 9 1 1 NMOS W=1u L=1u
R2 2 VDD 1k
M3 2 7 12 12 NMOS W=1u L=1u
R1 4 VDD 1k
M1 4 7 11 13 13 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

