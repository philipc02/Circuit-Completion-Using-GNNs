*SPICE Netlist for circuit 531
M1 5 1 0 12 12 NMOS W=1u L=1u
M4 3 1 0 0 NMOS W=1u L=1u
R2 2 VDD 1k
M2 2 9 3 3 NMOS W=1u L=1u
R3 5 3 1k
R1 4 VDD 1k
M3 4 8 5 5 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

