*SPICE Netlist for circuit 189
I1 1 0 DC 1mA
M2 2 7 1 1 NMOS W=1u L=1u
M1 3 5 1 1 NMOS W=1u L=1u
R1 2 VDD 1k
R2 3 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

