*SPICE Netlist for circuit 289
R3 0 3 1k
R2 3 1 1k
R1 1 VDD 1k
M1 1 5 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

