*SPICE Netlist for circuit 725
C1 2 VDD 1nF
C2 6 3 1nF
M2 6 1 2 2 PMOS W=1u L=1u
R1 0 3 1k
M1 3 2 VDD VDD PMOS W=1u L=1u
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

