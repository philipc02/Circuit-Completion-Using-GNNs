*SPICE Netlist for circuit 332
I1 VDD 4 DC 1mA
V1 6 0 5V
M2 4 4 0 0 NMOS W=1u L=1u
M3 3 4 0 0 NMOS W=1u L=1u
M1 6 3 4 4 NMOS W=1u L=1u
R1 3 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

