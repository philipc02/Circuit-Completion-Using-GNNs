*SPICE Netlist for circuit 557
C1 2 5 1nF
V1 5 0 5V
C2 0 2 1nF
I1 3 0 DC 1mA
R1 1 VDD 1k
M1 1 2 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

