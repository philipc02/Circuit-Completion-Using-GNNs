*SPICE Netlist for circuit 183
C1 3 4 1nF
M1 4 3 5 5 NMOS W=1u L=1u
M2 5 2 0 0 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

