*SPICE Netlist for circuit 751
C1 7 27 1nF
R2 27 3 1k
C2 8 28 1nF
R3 28 1 1k
R4 1 2 1k
R1 3 4 1k

.OP
.END

