*SPICE Netlist for circuit 369
C1 2 1 1nF
I1 2 0 DC 1mA
R1 3 1 1k
M1 VDD 1 2 2 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

