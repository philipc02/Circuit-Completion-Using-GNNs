*SPICE Netlist for circuit 703
C1 0 6 1nF
C2 0 3 1nF
M1 10 8 0 14 14 NMOS W=1u L=1u
M4 6 8 0 0 NMOS W=1u L=1u
M3 3 7 0 0 NMOS W=1u L=1u
M2 15 7 0 16 16 NMOS W=1u L=1u
M5 1 1 VDD VDD PMOS W=1u L=1u
M7 2 1 VDD VDD PMOS W=1u L=1u
M6 15 2 VDD VDD PMOS W=1u L=1u
M8 2 2 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

