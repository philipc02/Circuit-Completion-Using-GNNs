*SPICE Netlist for circuit 685
C1 2 1 1nF
R1 5 1 1k

.OP
.END

