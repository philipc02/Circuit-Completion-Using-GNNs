*SPICE Netlist for circuit 318
C1 3 2 1nF
M2 3 6 0 0 NMOS W=1u L=1u
M3 4 1 0 0 NMOS W=1u L=1u
M1 VDD 2 4 4 NMOS W=1u L=1u
R2 2 VDD 1k
R1 3 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

