*SPICE Netlist for circuit 749
R2 1 4 1k
R4 1 5 1k
R1 7 1 1k
R3 8 1 1k

.OP
.END

