*SPICE Netlist for circuit 284
V1 1 0 5V
R1 2 0 1k
M1 1 2 0 0 PMOS W=1u L=1u
R2 2 1 1k
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

