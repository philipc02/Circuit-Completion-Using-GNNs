*SPICE Netlist for circuit 560
C1 4 2 1nF
C2 0 4 1nF
V1 3 0 5V
M2 3 4 0 0 NMOS W=1u L=1u
M1 2 1 3 3 NMOS W=1u L=1u
R1 2 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

