*SPICE Netlist for circuit 422
C1 2 VDD 1nF
C2 16 7 1nF
R3 10 16 1k
I1 3 0 DC 1mA
M1 8 1 10 17 17 NMOS W=1u L=1u
M5 8 2 VDD VDD NMOS W=1u L=1u
M6 5 2 VDD VDD PMOS W=1u L=1u
M4 10 13 3 3 NMOS W=1u L=1u
M2 7 14 3 3 NMOS W=1u L=1u
R2 8 2 1k
R1 2 5 1k
M3 5 1 7 7 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

