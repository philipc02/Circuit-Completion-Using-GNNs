*SPICE Netlist for circuit 342
C1 0 4 1nF
M3 5 2 4 4 NMOS W=1u L=1u
I1 VDD 2 DC 1mA
M1 2 2 0 0 NMOS W=1u L=1u
M2 6 1 5 5 NMOS W=1u L=1u
R1 6 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

