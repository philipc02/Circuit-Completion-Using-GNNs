*SPICE Netlist for circuit 576
R2 0 3 1k
R3 0 1 1k
R4 3 1 1k
M2 1 2 VDD VDD PMOS W=1u L=1u
R1 2 VDD 1k
M1 2 5 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

