*SPICE Netlist for circuit 262
I1 VDD 3 DC 1mA
M2 4 4 0 0 NMOS W=1u L=1u
R1 1 3 1k
M1 1 3 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

