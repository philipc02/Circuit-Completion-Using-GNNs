*SPICE Netlist for circuit 200
M1 1 0 3 3 NMOS W=1u L=1u
V1 4 0 5V
R1 1 VDD 1k
R2 4 3 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

