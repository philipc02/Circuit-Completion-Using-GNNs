*SPICE Netlist for circuit 654
M3 6 3 0 0 NMOS W=1u L=1u
M4 4 8 0 0 NMOS W=1u L=1u
M5 6 4 0 0 NMOS W=1u L=1u
M6 10 1 VDD VDD PMOS W=1u L=1u
M2 7 2 6 6 NMOS W=1u L=1u
M1 9 7 4 4 NMOS W=1u L=1u
M7 7 5 10 10 PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

