*SPICE Netlist for circuit 98
M2 1 4 0 0 NMOS W=1u L=1u
R1 0 2 1k
M1 VDD 1 2 2 NMOS W=1u L=1u
R2 1 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

