*SPICE Netlist for circuit 438
I1 VDD 1 DC 1mA
I2 1 0 DC 1mA
M1 1 0 0 0 NMOS W=1u L=1u
R1 1 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

