*SPICE Netlist for circuit 639
R1 0 4 1k
M4 4 7 0 0 PMOS W=1u L=1u
M2 8 1 VDD VDD PMOS W=1u L=1u
M3 5 2 8 8 PMOS W=1u L=1u
M1 5 3 4 4 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

