*SPICE Netlist for circuit 238
M3 1 3 0 0 NMOS W=1u L=1u
M2 5 9 1 1 NMOS W=1u L=1u
M1 4 7 1 1 NMOS W=1u L=1u
M4 5 2 10 11 11 PMOS W=1u L=1u
M5 4 2 12 12 PMOS W=1u L=1u
R1 10 VDD 1k
R2 12 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

