*SPICE Netlist for circuit 534
I1 VDD 5 DC 1mA
I2 VDD 3 DC 1mA
I3 6 0 DC 1mA
I4 4 0 DC 1mA
R1 6 4 1k
M4 6 5 VDD VDD PMOS W=1u L=1u
M3 4 3 VDD VDD PMOS W=1u L=1u
M1 3 7 4 4 NMOS W=1u L=1u
M2 5 8 6 6 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

