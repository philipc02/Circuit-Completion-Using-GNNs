*SPICE Netlist for circuit 197
V1 5 0 5V
M1 1 0 6 6 NMOS W=1u L=1u
R1 1 VDD 1k
R2 2 VDD 1k
M2 2 5 6 6 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

