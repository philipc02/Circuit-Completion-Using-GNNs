*SPICE Netlist for circuit 322
M1 1 1 0 0 NMOS W=1u L=1u
M2 3 1 0 0 NMOS W=1u L=1u
R3 1 3 1k
R2 3 VDD 1k
R1 1 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

