*SPICE Netlist for circuit 36
V1 4 0 5V
R1 0 2 1k
M1 4 1 2 2 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

