*SPICE Netlist for circuit 177
M2 3 2 0 0 NMOS W=1u L=1u
M3 6 1 VDD VDD PMOS W=1u L=1u
M1 6 5 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

