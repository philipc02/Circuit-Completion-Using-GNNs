*SPICE Netlist for circuit 386
C1 0 3 1nF
C2 0 4 1nF
C3 1 0 1nF
R3 0 3 1k
R2 1 VDD 1k
M2 1 7 3 3 NMOS W=1u L=1u
M1 4 7 3 8 8 NMOS W=1u L=1u
R1 4 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

