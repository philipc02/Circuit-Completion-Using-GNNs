*SPICE Netlist for circuit 599
C1 0 1 1nF
M1 2 6 0 0 NMOS W=1u L=1u
M2 1 0 4 4 NMOS W=1u L=1u
V1 6 0 5V
R3 0 4 1k
R4 4 2 1k
R1 2 VDD 1k
R2 1 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

