*SPICE Netlist for circuit 249
M5 2 1 0 0 NMOS W=1u L=1u
M4 7 11 2 2 NMOS W=1u L=1u
M2 13 9 2 2 NMOS W=1u L=1u
M1 4 3 7 14 14 NMOS W=1u L=1u
R1 4 VDD 1k
R2 5 VDD 1k
R3 7 5 1k
M3 5 3 13 13 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

