*SPICE Netlist for circuit 600
C1 1 4 1nF
I1 4 0 DC 1mA
M1 1 0 5 5 NMOS W=1u L=1u
V1 7 0 5V
R2 0 5 1k
R4 5 4 1k
R1 4 VDD 1k
R3 1 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

