*SPICE Netlist for circuit 363
C1 0 1 1nF
C2 0 3 1nF
C3 3 1 1nF
M1 1 3 0 0 NMOS W=1u L=1u
R1 1 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

