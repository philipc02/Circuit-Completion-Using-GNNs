*SPICE Netlist for circuit 604
M2 3 2 0 0 NMOS W=1u L=1u
V1 5 0 5V
R2 0 1 1k
R4 2 1 1k
M1 VDD 3 1 1 NMOS W=1u L=1u
R3 5 2 1k
R1 3 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

