*SPICE Netlist for circuit 360
I1 3 0 DC 1mA
V1 5 0 5V
R1 1 VDD 1k
M1 1 2 3 3 NMOS W=1u L=1u
R2 5 3 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

