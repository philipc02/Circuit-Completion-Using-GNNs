*SPICE Netlist for circuit 529
M1 2 4 0 0 NMOS W=1u L=1u
M2 2 1 5 5 PMOS W=1u L=1u
R1 5 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

