*SPICE Netlist for circuit 306
C1 9 VDD 1nF
C2 7 1 1nF
I1 VDD 2 DC 1mA
M2 3 1 0 0 NMOS W=1u L=1u
M1 2 2 0 0 NMOS W=1u L=1u
R1 2 1 1k
R2 9 3 1k
M3 3 8 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

