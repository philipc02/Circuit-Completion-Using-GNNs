*SPICE Netlist for circuit 594
I1 VDD 1 DC 1mA
M1 2 0 1 1 NMOS W=1u L=1u
R2 0 1 1k
R1 2 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

