*SPICE Netlist for circuit 93
R2 0 1 1k
M1 3 0 1 1 NMOS W=1u L=1u
R1 2 1 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

