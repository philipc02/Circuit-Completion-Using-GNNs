*SPICE Netlist for circuit 564
I1 3 0 DC 1mA
R1 0 4 1k
M3 1 1 VDD VDD PMOS W=1u L=1u
M4 2 1 VDD VDD PMOS W=1u L=1u
R2 4 2 1k
M2 1 8 3 3 NMOS W=1u L=1u
M1 2 4 3 3 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

