*SPICE Netlist for circuit 309
M1 2 1 0 0 NMOS W=1u L=1u
R1 1 2 1k
M2 2 1 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

