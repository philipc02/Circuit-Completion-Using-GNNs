*SPICE Netlist for circuit 708
I1 4 0 DC 1mA
M5 12 1 VDD 13 13 PMOS W=1u L=1u
M6 6 2 12 14 14 PMOS W=1u L=1u
M1 6 3 15 16 16 NMOS W=1u L=1u
M4 15 9 4 4 NMOS W=1u L=1u
M2 17 10 4 4 NMOS W=1u L=1u
M8 5 2 18 18 PMOS W=1u L=1u
M3 5 3 17 17 NMOS W=1u L=1u
M7 18 1 VDD VDD PMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)
.MODEL PMOS PMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

