*SPICE Netlist for circuit 54
C1 1 2 1nF
V1 1 0 5V
M1 VDD 1 2 2 NMOS W=1u L=1u
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

