*SPICE Netlist for circuit 231
M3 3 9 1 1 NMOS W=1u L=1u
M1 4 12 1 1 NMOS W=1u L=1u
M4 4 10 2 2 NMOS W=1u L=1u
M2 6 11 2 2 NMOS W=1u L=1u
R1 3 VDD 1k
R2 6 VDD 1k
.MODEL NMOS NMOS (LEVEL=1 VTO=1 KP=1.0e-4 LAMBDA=0.02)

.OP
.END

